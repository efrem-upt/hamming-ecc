module mux_5s_1b (
  input [0:31] i,
  input [4:0] s,
  output reg o);
  
always @(*) begin
  case (s)
    5'b00000: o = i[0];
    5'b00001: o = i[1];
    5'b00010: o = i[2];
    5'b00011: o = i[3];
    5'b00100: o = i[4];
    5'b00101: o = i[5];
    5'b00110: o = i[6];
    5'b00111: o = i[7];
    5'b01000: o = i[8];
    5'b01001: o = i[9];
    5'b01010: o = i[10];
    5'b01011: o = i[11];
    5'b01100: o = i[12];
    5'b01101: o = i[13];
    5'b01110: o = i[14];
    5'b01111: o = i[15];
    5'b10000: o = i[16];
    5'b10001: o = i[17];
    5'b10010: o = i[18];
    5'b10011: o = i[19];
    5'b10100: o = i[20];
    5'b10101: o = i[21];
    5'b10110: o = i[22];
    5'b10111: o = i[23];
    5'b11000: o = i[24];
    5'b11001: o = i[25];
    5'b11010: o = i[26];
    5'b11011: o = i[27];
    5'b11100: o = i[28];
    5'b11101: o = i[29];
    5'b11110: o = i[30];
    5'b11111: o = i[31];
  endcase
end
endmodule